-- Pieter-Jan Steeman

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY correlator_rx_test IS
END correlator_rx_test;

ARCHITECTURE structural OF correlator_rx_test IS

COMPONENT correlator_rx  -- component declaratie
	PORT
	(
		clk          	: IN  std_logic;		-- klok
		clk_en       	: IN  std_logic;		-- klok enable om kloksnelheid te verminderen
		rst          	: IN  std_logic;		-- reset
		sdi_despread 	: IN  std_logic;
		bit_sample   	: IN  std_logic;
		chip_sample2 	: IN  std_logic;
		data_out	: OUT std_logic
	);
END COMPONENT;

FOR uut : correlator_rx USE ENTITY work.correlator_rx(behavior); -- signalen aanmaken die overeenkomen met de poorten
  
	CONSTANT period   	: TIME := 100 ns;
	CONSTANT delay    	: TIME := 10 ns;
	SIGNAL end_of_sim 	: BOOLEAN := false;
	
	SIGNAL clk        	: std_logic;
	SIGNAL clk_en     	: std_logic;
	SIGNAL rst        	: std_logic;
	SIGNAL sdi_despread 	: std_logic;
	SIGNAL bit_sample 	: std_logic;
	SIGNAL chip_sample2	: std_logic;
	SIGNAL data_out    	: std_logic;
	
BEGIN

uut: correlator_rx PORT MAP -- ports aan signalen verbinden met port mapping
    (
      	clk    	   		=> clk,
      	clk_en 		   	=> clk_en,
      	rst    		   	=> rst,
      	sdi_despread 		=> sdi_despread,
      	bit_sample 		=> bit_sample,
	chip_sample2		=> chip_sample2,
	data_out    		=> data_out
    );

clock : PROCESS -- kloksignaal aanmaken voor de synchrone elementen
	BEGIN
    	clk <= '0';
    	WAIT FOR period/2;
    	LOOP
			clk <= '0';
			WAIT FOR period/2;
			clk <= '1';
			WAIT FOR period/2;
			EXIT WHEN end_of_sim;
		END LOOP;
	WAIT;
  END PROCESS clock;

tb : PROCESS -- testbench

	PROCEDURE tbvector(CONSTANT stimvect : IN std_logic_vector(3 DOWNTO 0))IS -- test vector aanmaken
	BEGIN	
		chip_sample2 <= stimvect(3);
		bit_sample <= stimvect(2);
		sdi_despread <= stimvect(1);
		rst <= stimvect(0); -- inputs "linken" met de vector
		WAIT FOR period;

	END tbvector;
	BEGIN	-- verschillende mogelijke scenario's aflopen

		clk_en <= '1';

		tbvector("0001");
		WAIT FOR period*5;
		tbvector("0100");
		WAIT FOR period*5;
		FOR i IN 0 TO 30 LOOP
			tbvector("1010");
			tbvector("0010");
			WAIT FOR period*5;
		END LOOP;
		tbvector("0100");
		tbvector("0000");
		WAIT FOR period*5;
		FOR i IN 0 TO 30 LOOP
			tbvector("1000");
			tbvector("0000");
			WAIT FOR period*5;
		END LOOP;
		tbvector("0100");
		tbvector("0000");
		WAIT FOR period*5;
		FOR i IN 0 TO 10 LOOP
			tbvector("1010");
			tbvector("0010");
			WAIT FOR period*5;
		END LOOP;
		FOR i IN 0 TO 20 LOOP
			tbvector("1000");
			tbvector("0000");
			WAIT FOR period*5;
		END LOOP;
		tbvector("0100");
		tbvector("0000");
		WAIT FOR period*10;

		end_of_sim <= true;
		WAIT;

	END PROCESS;
END;



