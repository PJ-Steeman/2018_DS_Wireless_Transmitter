-- Pieter-Jan Steeman

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY shiftreg_rx_test IS
END shiftreg_rx_test;

ARCHITECTURE structural OF shiftreg_rx_test IS

COMPONENT shiftreg_rx  -- component declaratie
	PORT
	(
		clk        : IN std_logic;
		clk_en     : IN std_logic;
		rst        : IN std_logic;
		data_in    : IN std_logic;
		bit_sample : IN std_logic;
		pre	   : OUT std_logic_vector(6 DOWNTO 0); 
		latch      : OUT std_logic_vector(3 DOWNTO 0) 
	);
END COMPONENT;

FOR uut : shiftreg_rx USE ENTITY work.shiftreg_rx(behavior); -- signalen aanmaken die overeenkomen met de poorten
  
	CONSTANT period   	: TIME := 100 ns;
	CONSTANT delay    	: TIME := 10 ns;
	SIGNAL end_of_sim 	: BOOLEAN := false;
	
	SIGNAL clk        	: std_logic;
	SIGNAL clk_en     	: std_logic;
	SIGNAL rst        	: std_logic;
	SIGNAL data_in  	: std_logic;
	SIGNAL bit_sample 	: std_logic;
	SIGNAL pre		: std_logic_vector(6 DOWNTO 0);
	SIGNAL latch		: std_logic_vector(3 DOWNTO 0);
	
BEGIN

uut: shiftreg_rx PORT MAP -- ports aan signalen verbinden met port mapping
    (
      	clk    	   	=> clk,
      	clk_en 		=> clk_en,
      	rst    		=> rst,
      	data_in 	=> data_in,
      	bit_sample 	=> bit_sample,
	pre		=> pre,
	latch		=> latch
    );

clock : PROCESS -- kloksignaal aanmaken voor de synchrone elementen
	BEGIN
    	clk <= '0';
    	WAIT FOR period/2;
    	LOOP
			clk <= '0';
			WAIT FOR period/2;
			clk <= '1';
			WAIT FOR period/2;
			EXIT WHEN end_of_sim;
		END LOOP;
	WAIT;
  END PROCESS clock;

tb : PROCESS -- testbench

	PROCEDURE tbvector(CONSTANT stimvect : IN std_logic_vector(2 DOWNTO 0))IS -- test vector aanmaken
		BEGIN
		 
		data_in <= stimvect(2);
		bit_sample <= stimvect(1);
		rst <= stimvect(0); -- inputs "linken" met de vector
      
			WAIT FOR period;
	END tbvector;
	BEGIN	-- verschillende mogelijke scenario's aflopen

		clk_en <= '1';

		tbvector("001");
		WAIT FOR period;
		tbvector("100");
		WAIT FOR period;
		tbvector("110");
		WAIT FOR period;
		tbvector("100");
		WAIT FOR period*4;
		tbvector("010");
		WAIT FOR period*6;
		tbvector("100");
		WAIT FOR period*8;
		tbvector("010");
		WAIT FOR period*0;
      
		end_of_sim <= true;
		WAIT;

	END PROCESS;
END;

